// Universidade de Sao Paulo
// MBA em seguranca de dados
//
// Igor Machado
//
// Decision Tree

module memory (
   input          clk,
   input          rst,
	
   input  [7:0]   addr,
   output [31:0]  data
);

   localparam NODE = {  32'h2_0041_0_48, // N0  (2,  65,    1,  72)
                        32'h6_0001_0_3F, // N1  (6,  1,     2,  63)
                        32'h5_0026_0_35, // N2  (5,  38,    3,  53)
                        32'h1_0001_0_1E, // N3  (1,  1,     4,  30)
                        32'h7_0001_0_12, // N4  (7,  1,     5,  18)
                        32'h2_0029_0_11, // N5  (2,  41,    6,  17)
                        32'hD_01FB_0_08, // N6  (13, 507,   7,  8 )
                        32'hF_FFFF_F_FF, // N7             (ACCEPT)
                        32'hD_0514_0_10, // N8  (13, 1300,  9,  16)
                        32'hD_0401_0_0E, // N9  (13, 1025,  10, 14)
								
                        32'h0_E637_0_0D, // N10 (0,  58935, 11, 13)
                        32'h0_4E7C_0_0C, // N11 (0,  20092, 12, 12)
                        32'hF_FFFF_0_FF, // N12              (DROP)
                        32'h0_E639_7_0C, // N13 (0,  58937, 7,  12)
                        32'h8_0001_7_0F, // N14 (8,  1,     7,  15)
                        32'h3_0004_C_07, // N15 (3,  4,     12, 7 )
                        32'hD_0599_7_07, // N16 (13, 1433,  7,  7 )
                        32'hD_000D_7_07, // N17 (13, 13,    7,  7 )
                        32'hD_0209_0_14, // N18 (13, 521,   19, 20)								
                        32'hD_01FB_7_0C, // N19 (13, 507,   7,  12)
								
                        32'hD_FFF4_0_1C, // N20 (13, 65524, 21, 28)
                        32'h2_002A_0_19, // N21 (2,  42,    22, 25)
                        32'hD_0428_0_07, // N22 (13, 1064,  23, 7 )
                        32'h3_0002_0_07, // N23 (3,  2,     24, 7 )
                        32'h0_ED46_7_07, // N24 (0,  60742, 7,  7 )
                        32'hD_0402_0_07, // N25 (13, 1026,  26, 7 )
                        32'h3_0004_0_07, // N26 (3,  4,     27, 7 )
                        32'hD_03A5_7_0C, // N27 (13, 933,   7,  12)
                        32'h3_0004_0_07, // N28 (3,  4,     29, 7 )
                        32'h5_0016_C_07, // N29 (5,  22,    12, 7 )
								
                        32'hD_0001_0_2B, // N30 (13, 1,     31, 43)
                        32'h0_003C_0_24, // N31 (0,  60,    32, 36)
                        32'hA_0001_0_23, // N32 (10, 1,     33, 35)
                        32'h3_0001_C_22, // N33 (3,  1,     12, 34)
                        32'h3_0005_7_07, // N34 (3,  5,     7,  7 )
                        32'h7_0001_7_07, // N35 (7,  1,     7,  7 )
                        32'h0_976F_7_25, // N36 (0,  38767, 7,  37)
                        32'h0_97B9_C_26, // N37 (0,  38841, 12, 38)
                        32'h0_A1FB_0_28, // N38 (0,  41467, 39, 40)
                        32'h0_A144_7_0C, // N39 (0,  41284, 7,  12)
								
                        32'h0_ED26_0_2A, // N40 (0,  60710, 41, 42)
                        32'hA_0001_7_07, // N41 (10, 1,     7,  7 )
                        32'h0_ED9B_C_07, // N42 (0,  60827, 12, 7 )
                        32'h4_0013_0_33, // N43 (4,  19,    44, 51)
                        32'hD_7110_7_2D, // N44 (13, 28944, 7,  45)
                        32'hD_7150_0_2F, // N45 (13, 29008, 46, 47)
                        32'h0_6735_7_0C, // N46 (0,  26421, 7,  12)
                        32'h8_0001_0_32, // N47 (8,  1,     48, 50)
                        32'h0_C7C7_7_31, // N48 (0,  51143, 7,  49)
                        32'h0_C7D9_C_07, // N49 (0,  51161, 12, 7 )
								
                        32'h2_002E_7_0C, // N50 (2,  46,    7,  12)
                        32'hD_5514_7_34, // N51 (13, 21780, 7,  52)
                        32'hD_B576_C_07, // N52 (13, 46454, 12, 7 )
                        32'hD_3D85_7_36, // N53 (13, 15749, 7,  54)
                        32'hD_FC08_0_3E, // N54 (13, 64520, 55, 62)
                        32'h0_000B_7_38, // N55 (0,  11,    7,  56)
                        32'hD_4058_0_3A, // N56 (13, 16472, 57, 58)
                        32'h2_003E_7_0C, // N57 (2,  62,    7,  12)
                        32'hD_FA9D_7_3B, // N58 (13, 64157, 7,  59)
                        32'h0_D8E7_0_0C, // N59 (0,  55527, 60, 12)
								
                        32'h0_D854_0_0C, // N60 (0,  55380, 61, 12)
                        32'h0_C60C_C_0C, // N61 (0,  50700, 12, 12)
                        32'h7_0001_7_07, // N62 (7,  1,     7,  7 )
                        32'hD_0200_7_40, // N63 (13, 512,   7,  64)
                        32'h0_0002_7_41, // N64 (0,  2,     7,  65)
                        32'hD_4072_0_07, // N65 (13, 16498, 66, 7 )
                        32'h3_0004_0_07, // N66 (3,  4,     67, 7 )
                        32'hA_0001_C_44, // N67 (10, 1,     12, 68)
                        32'hD_0400_7_45, // N68 (13, 1024,  7,  69)
                        32'hD_3D00_0_0C, // N69 (13, 15616, 70, 12)
								
                        32'hD_0401_0_07, // N70 (13, 1025,  71, 7 )
                        32'h1_0001_C_07, // N71 (1,  1,     12, 7 )
                        32'h9_0001_7_07  // N72 (9,  1,     7,  7 )
                     };
							
   reg [31:0] data_mem;
   reg [31:0] data_mem_ff;

   always @(*)
   begin
      case(addr)
         8'h0:    data_mem = NODE[2335:2304];
         8'h1:    data_mem = NODE[2303:2272];
         8'h2:    data_mem = NODE[2271:2240]; 
         8'h3:    data_mem = NODE[2239:2208];
         8'h4:    data_mem = NODE[2207:2176];
         8'h5:    data_mem = NODE[2175:2144];
         8'h6:    data_mem = NODE[2143:2112];
         8'h7:    data_mem = NODE[2111:2080];
         8'h8:    data_mem = NODE[2079:2048];
         8'h9:    data_mem = NODE[2047:2016];
         8'hA:    data_mem = NODE[2015:1984];
         8'hB:    data_mem = NODE[1983:1952];
         8'hC:    data_mem = NODE[1951:1920];
         8'hD:    data_mem = NODE[1919:1888];
         8'hE:    data_mem = NODE[1887:1856];
         8'hF:    data_mem = NODE[1855:1824];
         8'h10:   data_mem = NODE[1823:1792];
         8'h11:   data_mem = NODE[1791:1760];
         8'h12:   data_mem = NODE[1759:1728];
         8'h13:   data_mem = NODE[1727:1696];
         8'h14:   data_mem = NODE[1695:1664];
         8'h15:   data_mem = NODE[1663:1632];
         8'h16:   data_mem = NODE[1631:1600];
         8'h17:   data_mem = NODE[1599:1568];
         8'h18:   data_mem = NODE[1567:1536];
         8'h19:   data_mem = NODE[1535:1504];
         8'h1A:   data_mem = NODE[1503:1472];
         8'h1B:   data_mem = NODE[1471:1440];
         8'h1C:   data_mem = NODE[1439:1408];
         8'h1D:   data_mem = NODE[1407:1376];
         8'h1E:   data_mem = NODE[1375:1344];
         8'h1F:   data_mem = NODE[1343:1312];
         8'h20:   data_mem = NODE[1311:1280];
         8'h21:   data_mem = NODE[1279:1248];
         8'h22:   data_mem = NODE[1247:1216];
         8'h23:   data_mem = NODE[1215:1184];
         8'h24:   data_mem = NODE[1183:1152];
         8'h25:   data_mem = NODE[1151:1120];
         8'h26:   data_mem = NODE[1119:1088];
         8'h27:   data_mem = NODE[1087:1056];
         8'h28:   data_mem = NODE[1055:1024];
         8'h29:   data_mem = NODE[1023:992];
         8'h2A:   data_mem = NODE[991:960];
         8'h2B:   data_mem = NODE[959:928];
         8'h2C:   data_mem = NODE[927:896];
         8'h2D:   data_mem = NODE[895:864];
         8'h2E:   data_mem = NODE[863:832];
         8'h2F:   data_mem = NODE[831:800];
         8'h30:   data_mem = NODE[799:768];
         8'h31:   data_mem = NODE[767:736];
         8'h32:   data_mem = NODE[735:704];
         8'h33:   data_mem = NODE[703:672];
         8'h34:   data_mem = NODE[671:640];
         8'h35:   data_mem = NODE[639:608];
         8'h36:   data_mem = NODE[607:576];
         8'h37:   data_mem = NODE[575:544];
         8'h38:   data_mem = NODE[543:512];
         8'h39:   data_mem = NODE[511:480];
         8'h3A:   data_mem = NODE[479:448];
         8'h3B:   data_mem = NODE[447:416];
         8'h3C:   data_mem = NODE[415:384];
         8'h3D:   data_mem = NODE[383:352];
         8'h3E:   data_mem = NODE[351:320];
         8'h3F:   data_mem = NODE[319:288];
         8'h40:   data_mem = NODE[287:256];
         8'h41:   data_mem = NODE[255:224];
         8'h42:   data_mem = NODE[223:192];
         8'h43:   data_mem = NODE[191:160];
         8'h44:   data_mem = NODE[159:128];
         8'h45:   data_mem = NODE[127:96];
         8'h46:   data_mem = NODE[95:64];
         8'h47:   data_mem = NODE[63:32];
         8'h48:   data_mem = NODE[31:0];
         default: data_mem = NODE[2335:2304];
   endcase
   end
	
   always @(posedge clk or posedge rst)
   begin
      if(rst)
      begin
         data_mem_ff <= NODE[2335:2304];
      end
		
      else
      begin
         data_mem_ff <= data_mem;
      end
   end
	
   assign data = data_mem_ff;
	
endmodule